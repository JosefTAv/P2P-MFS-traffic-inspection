../../../IPs/packet_detect/packet_detect.sv