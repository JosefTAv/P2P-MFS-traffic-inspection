../../../IPs/clk_sync_pulse/clk_sync_pulse.sv