../../../IPs/timestamp_inject/timestamp_inject.sv