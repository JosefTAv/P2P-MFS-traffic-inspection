../../../IPs/clk_sync_pulse/clk_sync_pulse_regs.sv